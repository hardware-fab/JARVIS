//`define IMPL_SOC
